******Sense_amplifier********


M00 gnd en   n1   gnd n w=1.8u l=0.4u
M01 n1  n2   nout gnd n w=1.8u l=0.4u
M02 n2  nout n1   gnd n w=1.8u l=0.4u
M03 vdd n2   nout vdd p w=3.6u l=0.4u
M04 n2  nout vdd  vdd p w=3.6u l=0.4u
M05 bl  en   nout vdd p w=4.8u l=0.4u
M06 n2  en   blb  vdd p w=4.8u l=0.4u
.END 

